--
--
--
--layers: for layer in 0 to N_LAYERS generate
--
--	for node in 0 to 
--
--end generate label;

library IEEE;
use IEEE.std_logic_1164.all;

library Work;
use Work.NetworkConstants.all;

entity NeuralNetwork is
	port(
		i_CLK: in std_logic
	);
end entity;

architecture nn of NeuralNetwork is
begin
	
end;
